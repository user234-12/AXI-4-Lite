class shared_container;
    static logic [31:0]shared_addr;
endclass
