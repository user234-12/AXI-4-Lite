`define WIDTH_ADDR 32
`define WIDTH_DATA 32
`define STROBE_WIDTH 32
`define NO_OF_SEQ 100
